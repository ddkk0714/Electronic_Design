module top(
    input clk,           // 100MHz �Է� Ŭ��
    input rst,
    input [7:0] btn,
    output piezo
);

    wire clk_1MHz;

    // Ŭ�� ����� ���
    clk_div_1MHz u_clk_div (
        .clk(clk),
        .rst(rst),
        .clk_1MHz(clk_1MHz)
    );

    // �ǿ��� ���
    piezo_basic u_piezo (
        .clk(clk_1MHz),
        .rst(rst),
        .btn(btn),
        .piezo(piezo)
    );

endmodule
