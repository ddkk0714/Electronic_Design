`timescale 1us/1ns

module tb_seg_counter;
reg clk;
reg rst;
reg btn;
wire [7:0] seg;

seg_counter UUT (
    .clk(clk),
    .rst(rst),
    .btn(btn),
    .seg(seg)
);

always begin
    #1 clk = ~clk; // 500kHz Ŭ��
end

initial begin
    clk = 0;
    rst = 1;
    btn = 0;

    // ����
    #10 rst = 0;
    #10 rst = 1;

    // ��ư ���� �׽�Ʈ
    #20 btn = 1;
    #10 btn = 0;
    
    #20 btn = 1;
    #10 btn = 0;

    #20 btn = 1;
    #10 btn = 0;
    
    #20 btn = 1;
    #10 btn = 0;
    
    #20 btn = 1;
    #10 btn = 0;
    
    #20 btn = 1;
    #10 btn = 0;
    
    #20 btn = 1;
    #10 btn = 0;
    
    #20 btn = 1;
    #10 btn = 0;
    
    #20 btn = 1;
    #10 btn = 0;
    
    #20 btn = 1;
    #10 btn = 0;
    
    #20 btn = 1;
    #10 btn = 0;
    #100 $finish;
end

endmodule
