`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/11/09 09:41:04
// Design Name: 
// Module Name: oneshot_universal
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module oneshot_universal #(
    parameter WIDTH = 1
)(
    input                  clk,
    input                  rst,             
    input  [WIDTH-1:0]     btn,              //���� ��Ʈ�� ����
    output reg [WIDTH-1:0] btn_trig
);
    // 2-FF ����ȭ
    reg [WIDTH-1:0] sync0, sync1;
    // ���� ���� ����(���� ���� ����)
    reg [WIDTH-1:0] prev;

    always @(posedge clk or negedge rst) begin
        if (!rst) begin
            sync0    <= {WIDTH{1'b0}};
            sync1    <= {WIDTH{1'b0}};
            prev     <= {WIDTH{1'b0}};
            btn_trig <= {WIDTH{1'b0}};
        end else begin
            sync0 <= btn;
            sync1 <= sync0;

            btn_trig <=  sync1 & ~prev;

            prev <= sync1;
        end
    end
endmodule

