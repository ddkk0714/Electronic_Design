module clk_div_1MHz(
    input clk,           // �Է�: 100MHz Ŭ��
    input rst,
    output reg clk_1MHz  // ���: 1MHz Ŭ��
);

    reg [7:0] cnt;  // 7��Ʈ�� 0~127 ���� (100���� ���)

    always @(posedge clk or negedge rst) begin
        if (!rst) begin
            cnt <= 0;
            clk_1MHz <= 0;
        end else if (cnt == 99) begin //1MHz�϶� 49, 5000KHz�϶� 99
            cnt <= 0;
            clk_1MHz <= ~clk_1MHz;  // 50 + 50 = 100 �� ���ֺ� 100
        end else begin
            cnt <= cnt + 1;
        end
    end
endmodule
